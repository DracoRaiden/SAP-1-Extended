module top_module;
    wire clk;
    ClockGenerator cg(clk);
endmodule